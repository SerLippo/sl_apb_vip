`ifndef APB_DEFINE_SV
`define APB_DEFINE_SV

`define ADDR_WIDTH 32
`define DATA_WIDTH 32

`endif