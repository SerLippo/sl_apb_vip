`ifndef APB_DEFINE_SV
`define APB_DEFINE_SV

`define ADDR_WIDTH 16
`define DATA_WIDTH 16

`endif