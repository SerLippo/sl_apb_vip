`ifndef APB_PKG_SV
`define APB_PKG_SV

`include "apb_define.sv"

package apb_test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import apb_pkg::*;

  `include "apb_env.sv"
  `include "apb_sequences.svh"
  `include "apb_tests.svh"

endpackage: apb_test_pkg

`endif