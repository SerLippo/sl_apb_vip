`ifndef APB_PKG_SV
`define APB_PKG_SV

`include "apb_define.sv"
`include "apb_if.sv"

package apb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_typedef.sv"
  `include "apb_config.sv"

  `include "apb_transaction.sv"
  `include "apb_master_seq_lib.sv"
  `include "apb_master_sequencer.sv"
  `include "apb_master_driver.sv"
  `include "apb_master_monitor.sv"
  `include "apb_master_agent.sv"
  `include "apb_slave_sequencer.sv"
  `include "apb_slave_driver.sv"
  `include "apb_slave_monitor.sv"
  `include "apb_slave_agent.sv"

endpackage: apb_pkg

`endif